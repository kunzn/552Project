
module CLA4 (
  input [3:0] A, 
  input [3:0] B, //Input values
  input Cin, // add-sub indicator
  output [3:0] Sum, //sum output
  output Ovfl, //To indicate overflow
  output Cout
);
	wire [3:0] carry;
	wire [3:0] p, g;
	wire [3:0] CoutTemp;

	assign g = A & B;
	assign p = A ^ B;

	assign carry[0] = Cin;
	assign carry[1] = g[0] | (p[0] & Cin); 
	assign carry[2] = g[1] | (p[1] & g[0]) | (p[1] & p[0] & Cin);
	assign carry[3] = g[2] | (p[2] & g[1]) | (p[2] & p[1] & g[0]) | (p[2] & p[1] & p[0] & Cin);
	assign Cout = g[3] | (p[3] & g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0]) | (p[3] & p[2] & p[1] & p[0] & Cin);

	assign Sum = p^carry;

	assign Ovfl = Cout ^ carry[3];
endmodule